// instruction memory
module IM(input  [8:2]  addr,output [31:0] outdata );

  reg  [31:0] ROM[127:0];
initial begin

ROM[0]=32'h20020005;
ROM[1]=32'h2003000c;
ROM[2]=32'h2067fff7;
ROM[3]=32'h2001004c;
ROM[4]=32'h0020f809;
ROM[5]=32'h00e22025;
ROM[6]=32'h00642824;
ROM[7]=32'h00a42820;
ROM[8]=32'h10a70017;
ROM[9]=32'h0064202a;
ROM[10]=32'h10800001;
ROM[11]=32'h20050000;
ROM[12]=32'h00e2202a;
ROM[13]=32'h00853820;
ROM[14]=32'h00e23822;
ROM[15]=32'hac670044;
ROM[16]=32'h8c020050;
ROM[17]=32'h08000020;
ROM[18]=32'h20020001;
ROM[19]=32'h00073840;
ROM[20]=32'h0c000017;
ROM[21]=32'h201f0014;
ROM[22]=32'h03e00008;
ROM[23]=32'h3c0155aa;
ROM[24]=32'h282155aa;
ROM[25]=32'h14200006;
ROM[26]=32'h34e70005;
ROM[27]=32'h30e10005;
ROM[28]=32'h00e10821;
ROM[29]=32'h00210823;
ROM[30]=32'h00073842;
ROM[31]=32'h03e00008;
ROM[32]=32'hac020054;
ROM[33]=32'h08000021;

/*
ROM[0]=32'h3c039876;
ROM[1]=32'h34021234;
ROM[2]=32'h00624023;
ROM[3]=32'h01034826;
ROM[4]=32'h01285021;
ROM[5]=32'h01425020;
ROM[6]=32'h01435822;
ROM[7]=32'h016a6027;
ROM[8]=32'h016a6825;
ROM[9]=32'h016a7024;
ROM[10]=32'h01ac982a;
ROM[11]=32'h01aca02b;
ROM[12]=32'h000840c0;
ROM[13]=32'h00084c02;
ROM[14]=32'h00085743;
ROM[15]=32'h340b3410;
ROM[16]=32'h01686004;
ROM[17]=32'h01686806;
ROM[18]=32'h01687007;
ROM[19]=32'h00432021;
ROM[20]=32'h201d0000;
ROM[21]=32'hafa40000;
ROM[22]=32'hafa40004;
ROM[23]=32'hafa40008;
ROM[24]=32'ha7a80004;
ROM[25]=32'ha7a9000a;
ROM[26]=32'ha3aa0007;
ROM[27]=32'ha3a80009;
ROM[28]=32'ha3a90008;
ROM[29]=32'h8fa80000;
ROM[30]=32'hafa8000c;
ROM[31]=32'h87a90002;
ROM[32]=32'hafa90010;
ROM[33]=32'h97a90002;
ROM[34]=32'hafa90014;
ROM[35]=32'h83aa0003;
ROM[36]=32'hafaa0018;
ROM[37]=32'h93aa0003;
ROM[38]=32'hafaa001c;
ROM[39]=32'h93aa0001;
ROM[40]=32'hafaa0020;
*/
/*
ROM[0]=32'h20020001;
ROM[1]=32'h20030001;
ROM[2]=32'h20070003;
ROM[3]=32'h00434020;
ROM[4]=32'h00031020;
ROM[5]=32'h00081820;
ROM[6]=32'h20e70001;
ROM[7]=32'h20e6fff6;
ROM[8]=32'h18c0fffa;
ROM[9]=32'h20020001;
ROM[10]=32'h20030001;
ROM[11]=32'h2007000a;
ROM[12]=32'h00434020;
ROM[13]=32'h00031020;
ROM[14]=32'h00081820;
ROM[15]=32'h20e7ffff;
ROM[16]=32'h20e6fffd;
ROM[17]=32'h04c1fffa;
ROM[18]=32'h20020001;
ROM[19]=32'h20030001;
ROM[20]=32'h2007000b;
ROM[21]=32'h00434020;
ROM[22]=32'h00031020;
ROM[23]=32'h00081820;
ROM[24]=32'h20e7ffff;
ROM[25]=32'h20e6fffd;
ROM[26]=32'h1cc0fffa;
ROM[27]=32'h20020001;
ROM[28]=32'h20030001;
ROM[29]=32'h20070003;
ROM[30]=32'h00434020;
ROM[31]=32'h00031020;
ROM[32]=32'h00081820;
ROM[33]=32'h20e70001;
ROM[34]=32'h20e6fff5;
ROM[35]=32'h04c0fffa;
ROM[36]=32'h2008ffff;
*/
/*
ROM[0]=32'h20020005;
ROM[1]=32'h2003000c;
ROM[2]=32'h2067fff7;
ROM[3]=32'h00e22025;
ROM[4]=32'h00642824;
ROM[5]=32'h00a42820;
ROM[6]=32'h10a7000a;
ROM[7]=32'h0064202a;
ROM[8]=32'h10800001;
ROM[9]=32'h20050000;
ROM[10]=32'h00e2202a;
ROM[11]=32'h00853820;
ROM[12]=32'h00e23822;
ROM[13]=32'hac670044;
ROM[14]=32'h8c020050;
ROM[15]=32'h08000011;
ROM[16]=32'h20020001;
ROM[17]=32'hac020054;
ROM[18]=32'h08000012;
*/
//$readmemh("C:\Users\lenovo3\Documents\Tencent Files\1756375671\FileRecv\test(2).txt", ROM);
end
  assign outdata = ROM[addr]; 
endmodule 
